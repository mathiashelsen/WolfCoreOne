-- This file contains all constant things, such as bit locations of the
-- instructions, addresses of IOs etc.

package mainArch is

constant IMM : natural := 31;
type REGA is range 30 downto 27;
type REGB is range 26 downto 23;

end package;
