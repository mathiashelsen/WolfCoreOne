library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity progMem is
	port(
		instrOutput	: out std_logic_vector(31 downto 0);
		instrAddress: in std_logic_vector(31 downto 0);
		clk			: in std_logic
	);
end entity;

architecture default of progMem is
	type regFileType is array(3 downto 0) of std_logic_vector(31 downto 0);
begin
process(clk) begin
	if (clk'event and clk='0') then
		case instrAddress is
			when X"0000_0004" =>
				instrOutput <= X"00000502";
			when X"0000_0005" =>
				instrOutput <= X"88002612";
			when X"0000_0006" =>
				instrOutput <= X"e80047d2";
			when others =>
				instrOutput <= X"0000_0000";
		end case;
	end if;
end process;
end architecture;
