library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package custom_types is
    type instruction is ( CLEAR, READOUT );
end custom_types;
